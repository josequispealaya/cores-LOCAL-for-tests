module And(
    input i_a,
    input i_b,
    output o_z
);

    assign o_z = i_a & i_b;

endmodule